** Profile: "SCHEMATIC1-Sim_Transient"  [ D:\FACULTATE\AN_1_MASTER\PAC\Teme\Tema5_EtajAmplClAB\tema5_etajamplclab-SCHEMATIC1-Sim_Transient.sim ] 

** Creating circuit file "tema5_etajamplclab-SCHEMATIC1-Sim_Transient.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tema5_etajamplclab-SCHEMATIC1.net" 


.END
